module test (
    
);
    reg i7,i6,i5,i4,i3,i2,i1,i0,s2,s1,s0;
    wire out;
    eightXoneMux a1(out,i7,i6,i5,i4,i3,i2,i1,i0,s2,s1,s0);
    initial begin
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 0;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 0;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 0;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 0;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 0;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 0;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 0;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 0;s2 = 1;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 0;s1 = 1;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 0;s0 = 1;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 0;#1
        i7 = 1;i6 = 1;i5 = 1;i4 = 1;i3 = 1;i2 = 1;i1 = 1;i0 = 1;s2 = 1;s1 = 1;s0 = 1;#1

        $finish;
    end
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0,a1);
    end
endmodule