`timescale 1ns/1ns
module test (
    
);
    reg i3,i2,i1,i0,s1,s0;
    wire out;
    fourXoneMux a1(out,i3,i2,i1,i0,s1,s0);
    initial begin
        i3=0;i2=0;i1=0;i0=0;s1=0;s0=0;#1
        i3=0;i2=0;i1=0;i0=0;s1=0;s0=1;#1
        i3=0;i2=0;i1=0;i0=0;s1=1;s0=0;#1
        i3=0;i2=0;i1=0;i0=0;s1=1;s0=1;#1
        i3=0;i2=0;i1=0;i0=1;s1=0;s0=0;#1
        i3=0;i2=0;i1=0;i0=1;s1=0;s0=1;#1
        i3=0;i2=0;i1=0;i0=1;s1=1;s0=0;#1
        i3=0;i2=0;i1=0;i0=1;s1=1;s0=1;#1
        i3=0;i2=0;i1=1;i0=0;s1=0;s0=0;#1
        i3=0;i2=0;i1=1;i0=0;s1=0;s0=1;#1
        i3=0;i2=0;i1=1;i0=0;s1=1;s0=0;#1
        i3=0;i2=0;i1=1;i0=0;s1=1;s0=1;#1
        i3=0;i2=0;i1=1;i0=1;s1=0;s0=0;#1
        i3=0;i2=0;i1=1;i0=1;s1=0;s0=1;#1
        i3=0;i2=0;i1=1;i0=1;s1=1;s0=0;#1
        i3=0;i2=0;i1=1;i0=1;s1=1;s0=1;#1
        i3=0;i2=1;i1=0;i0=0;s1=0;s0=0;#1
        i3=0;i2=1;i1=0;i0=0;s1=0;s0=1;#1
        i3=0;i2=1;i1=0;i0=0;s1=1;s0=0;#1
        i3=0;i2=1;i1=0;i0=0;s1=1;s0=1;#1
        i3=0;i2=1;i1=0;i0=1;s1=0;s0=0;#1
        i3=0;i2=1;i1=0;i0=1;s1=0;s0=1;#1
        i3=0;i2=1;i1=0;i0=1;s1=1;s0=0;#1
        i3=0;i2=1;i1=0;i0=1;s1=1;s0=1;#1
        i3=0;i2=1;i1=1;i0=0;s1=0;s0=0;#1
        i3=0;i2=1;i1=1;i0=0;s1=0;s0=1;#1
        i3=0;i2=1;i1=1;i0=0;s1=1;s0=0;#1
        i3=0;i2=1;i1=1;i0=0;s1=1;s0=1;#1
        i3=0;i2=1;i1=1;i0=1;s1=0;s0=0;#1
        i3=0;i2=1;i1=1;i0=1;s1=0;s0=1;#1
        i3=0;i2=1;i1=1;i0=1;s1=1;s0=0;#1
        i3=0;i2=1;i1=1;i0=1;s1=1;s0=1;#1
        i3=1;i2=0;i1=0;i0=0;s1=0;s0=0;#1
        i3=1;i2=0;i1=0;i0=0;s1=0;s0=1;#1
        i3=1;i2=0;i1=0;i0=0;s1=1;s0=0;#1
        i3=1;i2=0;i1=0;i0=0;s1=1;s0=1;#1
        i3=1;i2=0;i1=0;i0=1;s1=0;s0=0;#1
        i3=1;i2=0;i1=0;i0=1;s1=0;s0=1;#1
        i3=1;i2=0;i1=0;i0=1;s1=1;s0=0;#1
        i3=1;i2=0;i1=0;i0=1;s1=1;s0=1;#1
        i3=1;i2=0;i1=1;i0=0;s1=0;s0=0;#1
        i3=1;i2=0;i1=1;i0=0;s1=0;s0=1;#1
        i3=1;i2=0;i1=1;i0=0;s1=1;s0=0;#1
        i3=1;i2=0;i1=1;i0=0;s1=1;s0=1;#1
        i3=1;i2=0;i1=1;i0=1;s1=0;s0=0;#1
        i3=1;i2=0;i1=1;i0=1;s1=0;s0=1;#1
        i3=1;i2=0;i1=1;i0=1;s1=1;s0=0;#1
        i3=1;i2=0;i1=1;i0=1;s1=1;s0=1;#1
        i3=1;i2=1;i1=0;i0=0;s1=0;s0=0;#1
        i3=1;i2=1;i1=0;i0=0;s1=0;s0=1;#1
        i3=1;i2=1;i1=0;i0=0;s1=1;s0=0;#1
        i3=1;i2=1;i1=0;i0=0;s1=1;s0=1;#1
        i3=1;i2=1;i1=0;i0=1;s1=0;s0=0;#1
        i3=1;i2=1;i1=0;i0=1;s1=0;s0=1;#1
        i3=1;i2=1;i1=0;i0=1;s1=1;s0=0;#1
        i3=1;i2=1;i1=0;i0=1;s1=1;s0=1;#1
        i3=1;i2=1;i1=1;i0=0;s1=0;s0=0;#1
        i3=1;i2=1;i1=1;i0=0;s1=0;s0=1;#1
        i3=1;i2=1;i1=1;i0=0;s1=1;s0=0;#1
        i3=1;i2=1;i1=1;i0=0;s1=1;s0=1;#1
        i3=1;i2=1;i1=1;i0=1;s1=0;s0=0;#1
        i3=1;i2=1;i1=1;i0=1;s1=0;s0=1;#1
        i3=1;i2=1;i1=1;i0=1;s1=1;s0=0;#1
        i3=1;i2=1;i1=1;i0=1;s1=1;s0=1;#1
        $finish;
    end
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0,a1);
    end
endmodule